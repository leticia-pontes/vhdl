LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY TB_PORTA_AND IS
END TB_PORTA_AND;

ARCHITECTURE TB OF TB_PORTA_AND IS
	COMPONENT PORTA_AND IS
		PORT (E1, E2: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
				S: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
	END COMPONENT;
	
	SIGNAL E1, E2, S: STD_LOGIC_VECTOR(7 DOWNTO 0);
BEGIN
	DUT: PORTA_AND
	PORT MAP (E1 => E1,
				 E2 => E2,
				 S  => S);
				 
	SIMULATION: PROCESS
	BEGIN
		E1 <= (OTHERS => '0');
		E2 <= (OTHERS => '0');
		
		WAIT FOR 100 NS;
		
		E1 <= "00001111";
		E2 <= "00000111";
		
		WAIT FOR 100 NS;
		
		E1 <= "00001111";
		E2 <= "00001111";
		
		WAIT;
	END PROCESS;
END TB;