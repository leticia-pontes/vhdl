LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY RELOGIO IS
    PORT (
        CLK : IN STD_LOGIC;
        RST : IN STD_LOGIC;
        A, B, C, D, E, F, G : OUT STD_LOGIC_VECTOR(5 DOWNTO 0)  -- 6 dígitos (HHMMSS)
    );
END RELOGIO;

ARCHITECTURE STRUCTURE OF RELOGIO IS

    -- Sinais BCD
    SIGNAL SEC_U, SEC_D : STD_LOGIC_VECTOR(3 DOWNTO 0); -- Segundos
    SIGNAL MIN_U, MIN_D : STD_LOGIC_VECTOR(3 DOWNTO 0); -- Minutos
    SIGNAL HRS_U, HRS_D : STD_LOGIC_VECTOR(3 DOWNTO 0); -- Horas

    -- Sinais de CARRY
    SIGNAL CARRY_SU, CARRY_SD, CARRY_MU, CARRY_MD, CARRY_HU : STD_LOGIC;

    -- Sinais dos segmentos para cada dígito
    SIGNAL SA, SB, SC, SD, SE, SF, SG : STD_LOGIC_VECTOR(5 DOWNTO 0);

    COMPONENT CONTADOR_BCD
        PORT (
            CLK     : IN STD_LOGIC;
            RST     : IN STD_LOGIC;
            ENABLE  : IN STD_LOGIC;
            BCD_OUT : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
            CARRY   : OUT STD_LOGIC
        );
    END COMPONENT;

    COMPONENT DECODER_BCD
        PORT (
            ENTRADA : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
            A, B, C, D, E, F, G : OUT STD_LOGIC
        );
    END COMPONENT;

BEGIN

    -- SEGUNDOS
    U1: CONTADOR_BCD PORT MAP (CLK => CLK, RST => RST, ENABLE => '1', BCD_OUT => SEC_U, CARRY => CARRY_SU);
    U2: CONTADOR_BCD PORT MAP (CLK => CLK, RST => RST, ENABLE => CARRY_SU, BCD_OUT => SEC_D, CARRY => CARRY_SD);

    -- MINUTOS
    U3: CONTADOR_BCD PORT MAP (CLK => CLK, RST => RST, ENABLE => CARRY_SD, BCD_OUT => MIN_U, CARRY => CARRY_MU);
    U4: CONTADOR_BCD PORT MAP (CLK => CLK, RST => RST, ENABLE => CARRY_MU, BCD_OUT => MIN_D, CARRY => CARRY_MD);

    -- HORAS
    U5: CONTADOR_BCD PORT MAP (CLK => CLK, RST => RST, ENABLE => CARRY_MD, BCD_OUT => HRS_U, CARRY => CARRY_HU);
    U6: CONTADOR_BCD PORT MAP (CLK => CLK, RST => RST, ENABLE => CARRY_HU, BCD_OUT => HRS_D, CARRY => OPEN);

    -- DECODIFICADORES
    D0: DECODER_BCD PORT MAP (ENTRADA => SEC_U, A => SA(0), B => SB(0), C => SC(0), D => SD(0), E => SE(0), F => SF(0), G => SG(0));
    D1: DECODER_BCD PORT MAP (ENTRADA => SEC_D, A => SA(1), B => SB(1), C => SC(1), D => SD(1), E => SE(1), F => SF(1), G => SG(1));
    D2: DECODER_BCD PORT MAP (ENTRADA => MIN_U, A => SA(2), B => SB(2), C => SC(2), D => SD(2), E => SE(2), F => SF(2), G => SG(2));
    D3: DECODER_BCD PORT MAP (ENTRADA => MIN_D, A => SA(3), B => SB(3), C => SC(3), D => SD(3), E => SE(3), F => SF(3), G => SG(3));
    D4: DECODER_BCD PORT MAP (ENTRADA => HRS_U, A => SA(4), B => SB(4), C => SC(4), D => SD(4), E => SE(4), F => SF(4), G => SG(4));
    D5: DECODER_BCD PORT MAP (ENTRADA => HRS_D, A => SA(5), B => SB(5), C => SC(5), D => SD(5), E => SE(5), F => SF(5), G => SG(5));

    -- SAÍDAS
    A <= SA; B <= SB; C <= SC; D <= SD; E <= SE; F <= SF; G <= SG;

END STRUCTURE;
