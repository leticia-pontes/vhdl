LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY COMPLEMENTO_DE_1 IS
	PORT (E1: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			S: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END COMPLEMENTO_DE_1;

ARCHITECTURE COMPLEMENTO_DE_1_ARCH OF COMPLEMENTO_DE_1 IS
BEGIN
	S <= NOT E1;
END COMPLEMENTO_DE_1_ARCH;