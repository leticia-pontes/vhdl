LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY PORTA_AND IS
	PORT (E1, E2: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			S: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END PORTA_AND;

ARCHITECTURE PORTA_AND_ARCH OF PORTA_AND IS
BEGIN
	S <= E1 AND E2;
END PORTA_AND_ARCH;