LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY COMPARAR IS
	PORT (E1, E2: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			S: OUT STD_LOGIC_VECTOR(2 DOWNTO 0));
END COMPARAR;

ARCHITECTURE COMPARAR_ARCH OF COMPARAR IS
BEGIN
	PROCESS(E1, E2)
	BEGIN
		IF E1 > E2 THEN
			S <= "010";
		ELSIF E1 < E2 THEN
			S <= "001";
		ELSIF E1 = E2 THEN
			S <= "100";
		END IF;
	END PROCESS;
END COMPARAR_ARCH;