LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY REGISTRADOR8BITS IS
	PORT (CLK, RST: IN STD_LOGIC;
			DIN: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			DOUT: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END REGISTRADOR8BITS;

ARCHITECTURE REGISTRADOR8BITS_ARCH OF REGISTRADOR8BITS IS
SIGNAL DADO: STD_LOGIC_VECTOR(7 DOWNTO 0);
BEGIN
	PROCESS(CLK, RST)
	BEGIN
		IF RST = '1' THEN
			DOUT <= (OTHERS => '0');
			DADO <= (OTHERS => '0');
		ELSIF (CLK'EVENT AND CLK = '1') THEN
			DADO <= DIN;
			DOUT <= DADO;
		END IF;
	END PROCESS;
END REGISTRADOR8BITS_ARCH;