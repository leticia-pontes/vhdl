LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY PORTA_XOR IS
	PORT (E1, E2: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			S: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END PORTA_XOR;

ARCHITECTURE PORTA_XOR_ARCH OF PORTA_XOR IS
BEGIN
	S <= E1 XOR E2;
END PORTA_XOR_ARCH;