LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY INCREMENTAR IS
	PORT (E1: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			S: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END INCREMENTAR;

ARCHITECTURE INCREMENTAR_ARCH OF INCREMENTAR IS
BEGIN
	S <= E1 + 1;
END INCREMENTAR_ARCH;