LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY ULA_COM_COMPARADOR IS
	PORT (CLK, RST: IN STD_LOGIC;
			A, B: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			SEL: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
			S: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END ULA_COM_COMPARADOR;

ARCHITECTURE ULA_COM_COMPARADOR_ARCH OF ULA_COM_COMPARADOR IS

COMPONENT PORTA_AND IS
	PORT (E1, E2: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			S: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END COMPONENT;

COMPONENT PORTA_OR IS
	PORT (E1, E2: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			S: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END COMPONENT;

COMPONENT PORTA_XOR IS
	PORT (E1, E2: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			S: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END COMPONENT;

COMPONENT ADICIONAR IS
	PORT (E1, E2: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			S: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END COMPONENT;

COMPONENT SUBTRAIR IS
	PORT (E1, E2: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			S: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END COMPONENT;

COMPONENT INCREMENTAR IS
	PORT (E1: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			S: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END COMPONENT;

COMPONENT DECREMENTAR IS
	PORT (E1: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			S: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END COMPONENT;

COMPONENT MUX3X8 IS
	PORT (E1, E2, E3, E4, E5, E6, E7: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			SEL: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
			S: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END COMPONENT;

COMPONENT REGISTRADOR8BITS IS
	PORT (CLK, RST: IN STD_LOGIC;
			DIN: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			DOUT: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END COMPONENT;

SIGNAL SIGNAL_A, SIGNAL_B, 
	RESULTADO_PORTA_AND, RESULTADO_PORTA_OR, RESULTADO_PORTA_XOR, 
	RESULTADO_ADICIONAR, RESULTADO_SUBTRAIR, RESULTADO_INCREMENTAR, RESULTADO_DECREMENTAR,
	RESULTADO_MUX3X8, RESULTADO_REGISTRADOR8BITS: STD_LOGIC_VECTOR(7 DOWNTO 0);

BEGIN
	-- REGISTRADORES
	REG_A: REGISTRADOR8BITS PORT MAP (CLK, RST, A, SIGNAL_A);
	REG_B: REGISTRADOR8BITS PORT MAP (CLK, RST, B, SIGNAL_B);

	-- OPERAÇÕES COM PORTAS
	OPERACAO_AND: PORTA_AND PORT MAP (SIGNAL_A, SIGNAL_B, RESULTADO_PORTA_AND);
	OPERACAO_OR: PORTA_OR PORT MAP (SIGNAL_A, SIGNAL_B, RESULTADO_PORTA_OR);
	OPERACAO_XOR: PORTA_XOR PORT MAP (SIGNAL_A, SIGNAL_B, RESULTADO_PORTA_XOR);
	
	-- OPERAÇÕES ARITMÉTICAS
	ADICAO: ADICIONAR PORT MAP (SIGNAL_A, SIGNAL_B, RESULTADO_ADICIONAR);
	SUBTRACAO: SUBTRAIR PORT MAP (SIGNAL_A, SIGNAL_B, RESULTADO_SUBTRAIR);
	
	-- OPERAÇÕES DE CONTAGEM
	INCREMENTO: INCREMENTAR PORT MAP (SIGNAL_A, RESULTADO_INCREMENTAR);
	DECREMENTO: DECREMENTAR PORT MAP (SIGNAL_A, RESULTADO_DECREMENTAR);
	
	-- MULTIPLEXADOR
	MUX: MUX3X8 PORT MAP (RESULTADO_PORTA_AND, RESULTADO_PORTA_OR, RESULTADO_PORTA_XOR, 
								 RESULTADO_ADICIONAR, RESULTADO_SUBTRAIR, RESULTADO_INCREMENTAR, RESULTADO_DECREMENTAR, 
								 SEL, RESULTADO_MUX3X8);
	
	REG3X8: REGISTRADOR8BITS PORT MAP (CLK, RST, RESULTADO_MUX3X8, S);
END ULA_COM_COMPARADOR_ARCH;






