LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY MULTIPLICAR_POR_2 IS
	PORT (E1: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			CARRY: OUT STD_LOGIC;
			S: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END MULTIPLICAR_POR_2;

ARCHITECTURE MULTIPLICAR_POR_2_ARCH OF MULTIPLICAR_POR_2 IS
BEGIN
	-- ATRIBUI O PRIMEIRO BIT AO CARRY
	CARRY <= E1(7);
	-- CONCATENA O RESTO DA ENTRADA COM O '0'
	S <= E1(6 DOWNTO 0) & '0';
END MULTIPLICAR_POR_2_ARCH;