LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY CONTADOR4BITS IS
	PORT(
		CLK, RST: IN STD_LOGIC;
		S: OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END CONTADOR4BITS;

ARCHITECTURE CONTADOR4BITS_ARCH OF CONTADOR4BITS IS
BEGIN
	PROCESS(CLK, RST)
	VARIABLE COUNT: STD_LOGIC_VECTOR(4 DOWNTO 0);
	BEGIN
		-- SE O RESET FOR ATIVADO
		IF RST = '1' THEN
			-- ZERA AS VARIÁVEIS
			COUNT := (OTHERS => '0'); -- CONTADOR
			S <= (OTHERS => '0'); -- SAÍDA
		-- SE FOR AÇÃO DO CLOCK (BORDA DE SUBIDA)
		ELSIF (CLK'EVENT AND CLK = '1') THEN
			-- SE FOR IGUAL A 16 (10000, 5 BITS)
			IF COUNT = "10000" THEN
				-- ZERA O CONTADOR
				COUNT := (OTHERS => '0');
			ELSE
				-- ATRIBUI O CONTADOR À SAÍDA, NO FORMATO 0000 (4 BITS)
				S <= COUNT(3 DOWNTO 0);
				-- INCREMENTA O CONTADOR
				COUNT := COUNT + 1;
			END IF;
		END IF;
	END PROCESS;
END CONTADOR4BITS_ARCH;
