LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY RELOGIO IS
    PORT (
        CLK_1HZ : IN STD_LOGIC;
        RST     : IN STD_LOGIC;
        -- SAÍDAS PARA OS 6 DÍGITOS
        SEG0_A, SEG0_B, SEG0_C, SEG0_D, SEG0_E, SEG0_F, SEG0_G : OUT STD_LOGIC;
        SEG1_A, SEG1_B, SEG1_C, SEG1_D, SEG1_E, SEG1_F, SEG1_G : OUT STD_LOGIC;
        SEG2_A, SEG2_B, SEG2_C, SEG2_D, SEG2_E, SEG2_F, SEG2_G : OUT STD_LOGIC;
        SEG3_A, SEG3_B, SEG3_C, SEG3_D, SEG3_E, SEG3_F, SEG3_G : OUT STD_LOGIC;
        SEG4_A, SEG4_B, SEG4_C, SEG4_D, SEG4_E, SEG4_F, SEG4_G : OUT STD_LOGIC;
        SEG5_A, SEG5_B, SEG5_C, SEG5_D, SEG5_E, SEG5_F, SEG5_G : OUT STD_LOGIC
    );
END RELOGIO;

ARCHITECTURE STRUCT OF RELOGIO IS
    COMPONENT CONT_BCD
        PORT (
            CLK     : IN STD_LOGIC;
            RST     : IN STD_LOGIC;
            ENABLE  : IN STD_LOGIC;
            BCD_OUT : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
            CARRY   : OUT STD_LOGIC
        );
    END COMPONENT;

    COMPONENT DECODER_BCD
        PORT (
            ENTRADA : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
            A, B, C, D, E, F, G : OUT STD_LOGIC
        );
    END COMPONENT;

    SIGNAL ENA : STD_LOGIC_VECTOR(5 DOWNTO 0); -- ENABLE
    SIGNAL CARRY : STD_LOGIC_VECTOR(5 DOWNTO 0);
    SIGNAL BCD : STD_LOGIC_VECTOR(3 DOWNTO 0) VECTOR(5 DOWNTO 0);
BEGIN
    -- PRIMEIRO CONTADOR (UNIDADE DE SEGUNDO)
    U0: CONT_BCD PORT MAP(CLK_1HZ, RST, '1', BCD(0), CARRY(0));
    -- DEMAIS CONTADORES COM ENTRADA DE CLOCK CONTROLADA PELO CARRY ANTERIOR
    U1: CONT_BCD PORT MAP(CLK_1HZ, RST, CARRY(0), BCD(1), CARRY(1));
    U2: CONT_BCD PORT MAP(CLK_1HZ, RST, CARRY(1), BCD(2), CARRY(2));
    U3: CONT_BCD PORT MAP(CLK_1HZ, RST, CARRY(2), BCD(3), CARRY(3));
    U4: CONT_BCD PORT MAP(CLK_1HZ, RST, CARRY(3), BCD(4), CARRY(4));
    U5: CONT_BCD PORT MAP(CLK_1HZ, RST, CARRY(4), BCD(5), CARRY(5));

    -- DECODIFICADORES
    D0: DECODER_BCD PORT MAP(BCD(0), SEG0_A, SEG0_B, SEG0_C, SEG0_D, SEG0_E, SEG0_F, SEG0_G);
    D1: DECODER_BCD PORT MAP(BCD(1), SEG1_A, SEG1_B, SEG1_C, SEG1_D, SEG1_E, SEG1_F, SEG1_G);
    D2: DECODER_BCD PORT MAP(BCD(2), SEG2_A, SEG2_B, SEG2_C, SEG2_D, SEG2_E, SEG2_F, SEG2_G);
    D3: DECODER_BCD PORT MAP(BCD(3), SEG3_A, SEG3_B, SEG3_C, SEG3_D, SEG3_E, SEG3_F, SEG3_G);
    D4: DECODER_BCD PORT MAP(BCD(4), SEG4_A, SEG4_B, SEG4_C, SEG4_D, SEG4_E, SEG4_F, SEG4_G);
    D5: DECODER_BCD PORT MAP(BCD(5), SEG5_A, SEG5_B, SEG5_C, SEG5_D, SEG5_E, SEG5_F, SEG5_G);
END STRUCT;
