LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY MUX2X4 IS
	PORT (E1, E2, E3, E4: IN STD_LOGIC;
			SEL: IN STD_LOGIC_VECTOR(1 DOWNTO 0);
			S: OUT STD_LOGIC);
END MUX2X4;

ARCHITECTURE MUX2X4_ARCH OF MUX2X4 IS
BEGIN
	PROCESS(SEL, E1, E2, E3, E4)
	BEGIN
		CASE SEL IS
			WHEN "00" => S <= E1;
			WHEN "01" => S <= E2;
			WHEN "10" => S <= E3;
			WHEN "11" => S <= E4;
			WHEN OTHERS => NULL;
		END CASE;
	END PROCESS;
END MUX2X4_ARCH;
