LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY COMPLEMENTO_DE_2 IS
	PORT (E1: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			S: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END COMPLEMENTO_DE_2;

ARCHITECTURE COMPLEMENTO_DE_2_ARCH OF COMPLEMENTO_DE_2 IS
BEGIN
	S <= (NOT E1) + 1;
END COMPLEMENTO_DE_2_ARCH;