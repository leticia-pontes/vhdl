LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY CONTADOR4BITS IS
	PORT(
		CLK, RST: IN STD_LOGIC;
		S: OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END CONTADOR4BITS;

ARCHITECTURE CONTADOR4BITS_ARCH OF CONTADOR4BITS IS
BEGIN
	PROCESS(CLK, RST)
	VARIABLE COUNT: STD_LOGIC_VECTOR(4 DOWNTO 0);
	BEGIN
		IF RST = '1' THEN
			-- ZERA AS VARIÁVEIS
			COUNT := (OTHERS => '0');
			S <= (OTHERS => '0');
		ELSIF (CLK'EVENT AND CLK = '1') THEN
			IF COUNT = "10000" THEN
				COUNT := (OTHERS => '0');
			ELSE
				S <= COUNT(3 DOWNTO 0);
				COUNT := COUNT + 1;
			END IF;
		END IF;
	END PROCESS;
END CONTADOR4BITS_ARCH;