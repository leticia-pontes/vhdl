LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY ULA IS
	PORT (CLK, RST: IN STD_LOGIC;
			A, B: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			SEL1, SEL2: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
			SEL_CARRY: IN STD_LOGIC_VECTOR(1 DOWNTO 0);
			MAIOR, MENOR, IGUAL, CARRY: OUT STD_LOGIC;
			S1, S2: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END ULA;

ARCHITECTURE ULA_ARCH OF ULA IS

COMPONENT PORTA_AND IS
	PORT (E1, E2: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			S: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END COMPONENT;

COMPONENT PORTA_OR IS
	PORT (E1, E2: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			S: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END COMPONENT;

COMPONENT PORTA_XOR IS
	PORT (E1, E2: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			S: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END COMPONENT;

COMPONENT ADICIONAR IS
	PORT (E1, E2: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			S: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END COMPONENT;

COMPONENT SUBTRAIR IS
	PORT (E1, E2: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			S: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END COMPONENT;

COMPONENT INCREMENTAR IS
	PORT (E1: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			S: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END COMPONENT;

COMPONENT DECREMENTAR IS
	PORT (E1: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			S: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END COMPONENT;

COMPONENT MUX3X8 IS
	PORT (E1, E2, E3, E4, E5, E6, E7: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			SEL: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
			S: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END COMPONENT;

COMPONENT REGISTRADOR8BITS IS
	PORT (CLK, RST: IN STD_LOGIC;
			DIN: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			DOUT: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END COMPONENT;

COMPONENT COMPARAR IS
	PORT (E1, E2: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			S: OUT STD_LOGIC_VECTOR(2 DOWNTO 0));
END COMPONENT;

COMPONENT DIVIDIR_POR_2 IS
	PORT (E1: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			CARRY: OUT STD_LOGIC;
			S: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END COMPONENT;

COMPONENT MULTIPLICAR_POR_2 IS
	PORT (E1: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			CARRY: OUT STD_LOGIC;
			S: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END COMPONENT;

COMPONENT COMPLEMENTO_DE_1 IS
	PORT (E1: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			S: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END COMPONENT;

COMPONENT COMPLEMENTO_DE_2 IS
	PORT (E1: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			S: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END COMPONENT;

COMPONENT MUX2X4 IS
	PORT (E1, E2, E3, E4: IN STD_LOGIC;
			SEL: IN STD_LOGIC_VECTOR(1 DOWNTO 0);
			S: OUT STD_LOGIC);
END COMPONENT;

SIGNAL SIGNAL_A, SIGNAL_B, 
	RESULTADO_PORTA_AND, RESULTADO_PORTA_OR, RESULTADO_PORTA_XOR, 
	RESULTADO_ADICIONAR, RESULTADO_SUBTRAIR, RESULTADO_INCREMENTAR, RESULTADO_DECREMENTAR,
	RESULTADO_MUX1, RESULTADO_MUX2, RESULTADO_REGISTRADOR8BITS, 
	RESULTADO_DIVIDIR, RESULTADO_MULTIPLICAR, 
	RESULTADO_COMPLEMENTO_DE_1, RESULTADO_COMPLEMENTO_DE_2: STD_LOGIC_VECTOR(7 DOWNTO 0);
	
SIGNAL RESULTADO_COMPARAR: STD_LOGIC_VECTOR(2 DOWNTO 0);

SIGNAL CARRY_DIVIDIR, CARRY_MULTIPLICAR, CARRY_FINAL: STD_LOGIC;

BEGIN
	-- REGISTRADORES
	REG_A: REGISTRADOR8BITS PORT MAP (CLK, RST, A, SIGNAL_A);
	REG_B: REGISTRADOR8BITS PORT MAP (CLK, RST, B, SIGNAL_B);

	-- OPERAÇÕES COM PORTAS
	OPERACAO_AND: PORTA_AND PORT MAP (SIGNAL_A, SIGNAL_B, RESULTADO_PORTA_AND);
	OPERACAO_OR: PORTA_OR PORT MAP (SIGNAL_A, SIGNAL_B, RESULTADO_PORTA_OR);
	OPERACAO_XOR: PORTA_XOR PORT MAP (SIGNAL_A, SIGNAL_B, RESULTADO_PORTA_XOR);
	
	-- OPERAÇÕES ARITMÉTICAS
	ADICAO: ADICIONAR PORT MAP (SIGNAL_A, SIGNAL_B, RESULTADO_ADICIONAR);
	SUBTRACAO: SUBTRAIR PORT MAP (SIGNAL_A, SIGNAL_B, RESULTADO_SUBTRAIR);
	
	-- OPERAÇÕES DE CONTAGEM
	INCREMENTO: INCREMENTAR PORT MAP (SIGNAL_A, RESULTADO_INCREMENTAR);
	DECREMENTO: DECREMENTAR PORT MAP (SIGNAL_A, RESULTADO_DECREMENTAR);
	
	-- MULTIPLEXADOR
	MUX1_3X8: MUX3X8 PORT MAP (RESULTADO_PORTA_AND, RESULTADO_PORTA_OR, RESULTADO_PORTA_XOR, 
										RESULTADO_ADICIONAR, RESULTADO_SUBTRAIR, RESULTADO_INCREMENTAR, RESULTADO_DECREMENTAR, 
										SEL1, RESULTADO_MUX1);
	
	-- REGISTRADOR DE 8 BITS
	REG_R1: REGISTRADOR8BITS PORT MAP (CLK, RST, RESULTADO_MUX1, S1);
	
	-- COMPARADOR
	COMPARACAO: COMPARAR PORT MAP(SIGNAL_A, SIGNAL_B, RESULTADO_COMPARAR);
	
	-- MULTIPLICAÇÃO E DIVISÃO POR 2
	DIVISAO: DIVIDIR_POR_2 PORT MAP(SIGNAL_A, CARRY_DIVIDIR, RESULTADO_DIVIDIR);
	MULTIPLICACAO: MULTIPLICAR_POR_2 PORT MAP(SIGNAL_A, CARRY_MULTIPLICAR, RESULTADO_MULTIPLICAR);
	
	-- COMPLEMENTOS DE 1 E 2
	OPERACAO_COMPLEMENTO_DE_1: COMPLEMENTO_DE_1 PORT MAP(SIGNAL_A, RESULTADO_COMPLEMENTO_DE_1);
	OPERACAO_COMPLEMENTO_DE_2: COMPLEMENTO_DE_2 PORT MAP(SIGNAL_A, RESULTADO_COMPLEMENTO_DE_2);
	
	-- MULTIPLEXADORES E REGISTRADORES
	MUX2_3X8: MUX3X8 PORT MAP (RESULTADO_MULTIPLICAR, RESULTADO_DIVIDIR, 
										RESULTADO_COMPLEMENTO_DE_1, RESULTADO_COMPLEMENTO_DE_2, 
										(OTHERS => '0'), (OTHERS => '0'), (OTHERS => '0'), 
										SEL2, RESULTADO_MUX2);
									
	-- REGISTRADOR DE 8 BITS
	REG_R2: REGISTRADOR8BITS PORT MAP (CLK, RST, RESULTADO_MUX2, S2);
	
	-- MULTIPLEXADOR
	MUX_2X4: MUX2X4 PORT MAP(CARRY_MULTIPLICAR, CARRY_DIVIDIR, '0', '0', SEL_CARRY, CARRY_FINAL);
	
	-- RESULTADOS
	MAIOR <= RESULTADO_COMPARAR(2);
	MENOR <= RESULTADO_COMPARAR(1);
	IGUAL <= RESULTADO_COMPARAR(0);
	CARRY <= CARRY_FINAL;
	
END ULA_ARCH;






