LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY ADICIONAR IS
	PORT (E1, E2: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			S: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END ADICIONAR;

ARCHITECTURE ADICIONAR_ARCH OF ADICIONAR IS
BEGIN
	S <= E1 + E2;
END ADICIONAR_ARCH;