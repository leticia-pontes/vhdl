LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY TB_DECODE3X8 IS
END TB_DECODE3X8;

ARCHITECTURE TB OF TB_DECODE3X8 IS
	COMPONENT DECODE3X8 IS
		PORT(
			CLK: IN STD_LOGIC;
			DIN: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
			DOUT: OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
		);
	END COMPONENT;
	
	SIGNAL CLK, PAUSE: STD_LOGIC;
	SIGNAL DIN: STD_LOGIC_VECTOR(2 DOWNTO 0);
	SIGNAL DOUT: STD_LOGIC_VECTOR(7 DOWNTO 0);
BEGIN
	DUT: DECODE3X8
		PORT MAP(CLK  => CLK,
					DIN  => DIN,
					DOUT => DOUT);
					
	CLK <= NOT CLK AFTER 50 NS WHEN PAUSE = '0' ELSE '0';
		
	STIMULI: PROCESS
	BEGIN
		PAUSE <= '0';
		
		DIN <= (OTHERS => '0');
		WAIT FOR 100 NS;
		
		DIN <= "001";
		WAIT FOR 100 NS;
		
		DIN <= "010";
		WAIT FOR 100 NS;
		
		DIN <= "011";
		WAIT FOR 100 NS;
		
		DIN <= "100";
		WAIT FOR 100 NS;
		
		DIN <= "101";
		WAIT FOR 100 NS;
		
		DIN <= "110";
		WAIT FOR 100 NS;
		
		DIN <= "111";
		WAIT FOR 100 NS;
		
		PAUSE <= '1';
		WAIT;
	END PROCESS;
END TB;