LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY DECREMENTAR IS
	PORT (E1: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			S: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END DECREMENTAR;

ARCHITECTURE DECREMENTAR_ARCH OF DECREMENTAR IS
BEGIN
	S <= E1 - 1;
END DECREMENTAR_ARCH;