LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY TB_RAM IS
END TB_RAM;

ARCHITECTURE TB OF TB_RAM IS
	-- COMPONENTE DA RAM
	COMPONENT RAM IS
		PORT(
			-- CLOCK, RESET, GRAVAÇÃO
			CLK, RST, WRITE_RAM: IN STD_LOGIC;
			-- ENDEREÇO DE DADO
			RAM_ADDR: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
			-- ENTRADA DE DADO
			RAM_DATAIN: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			-- SAÍDA DE DADO
			RAM_DATAOUT: OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
		);
	END COMPONENT;
	
	SIGNAL CLK, RST, WRITE_RAM, PAUSE: STD_LOGIC;
	SIGNAL RAM_DATAIN, RAM_DATAOUT: STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL RAM_ADDR: STD_LOGIC_VECTOR(4 DOWNTO 0);
BEGIN
	DUT: RAM
		PORT MAP (
			CLK => CLK,
			RST => RST,
			WRITE_RAM => WRITE_RAM,
			RAM_ADDR => RAM_ADDR,
			RAM_DATAIN => RAM_DATAIN,
			RAM_DATAOUT => RAM_DATAOUT
		);
		
	CLK <= NOT CLK AFTER 50 NS WHEN PAUSE = '0' ELSE '0';
	
	STIMULI: PROCESS
	BEGIN
		PAUSE <= '0';
		
		RST <= '0';
		WRITE_RAM <= '0';
		RAM_ADDR <= (OTHERS => '0');
		RAM_DATAIN <= (OTHERS => '0');
		WAIT FOR 100 NS;
		
		RAM_ADDR <= "00000";
		RAM_DATAIN <= "00000101";
		WRITE_RAM <= '1';
		WAIT FOR 100 NS;
		
		WRITE_RAM <= '0';
		WAIT FOR 100 NS;
		
		RAM_ADDR <= "00001";
		RAM_DATAIN <= "00001010";
		WRITE_RAM <= '1';
		WAIT FOR 100 NS;
		
		WRITE_RAM <= '0';
		WAIT FOR 100 NS;
		
		RAM_ADDR <= "00010";
		RAM_DATAIN <= "00001111";
		WRITE_RAM <= '1';
		WAIT FOR 100 NS;
		
		WRITE_RAM <= '0';
		WAIT FOR 100 NS;
		
		RAM_ADDR <= "01000";
		RAM_DATAIN <= "11111111";
		WRITE_RAM <= '1';
		WAIT FOR 100 NS;
		
		WRITE_RAM <= '0';
		WAIT FOR 100 NS;
		
		RAM_ADDR <= "00000";
		WAIT FOR 100 NS;
		
		RAM_ADDR <= "00001";
		WAIT FOR 100 NS;
		
		RAM_ADDR <= "00010";
		WAIT FOR 100 NS;
		
		RAM_ADDR <= "01000";
		WAIT FOR 100 NS;
		
		WAIT FOR 2000 NS;
		PAUSE <= '1';
		
		WAIT;
	END PROCESS;
END TB;