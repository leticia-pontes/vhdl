LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY PORTA_OR IS
	PORT (E1, E2: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			S: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END PORTA_OR;

ARCHITECTURE PORTA_OR_ARCH OF PORTA_OR IS
BEGIN
	S <= E1 OR E2;
END PORTA_OR_ARCH;