LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY CONTADOR4BITS IS
	PORT(
		CLK, RST, LOAD: IN STD_LOGIC;
		DIN: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		S: OUT STD_LOGIC_VECTOR(4 DOWNTO 0)
	);
END CONTADOR4BITS;

ARCHITECTURE CONTADOR4BITS_ARCH OF CONTADOR4BITS IS
BEGIN
	PROCESS(CLK, RST)
	VARIABLE COUNT: STD_LOGIC_VECTOR(4 DOWNTO 0);
	BEGIN
		-- SE O RESET FOR ATIVADO
		IF RST = '1' THEN
			-- ZERA AS VARIÁVEIS
			COUNT := (OTHERS => '0'); -- CONTADOR
			S <= (OTHERS => '0'); -- SAÍDA
		-- SE FOR AÇÃO DO CONTADOR
		ELSIF (CLK'EVENT AND CLK = '1') THEN
			-- SE FOR IGUAL A 16
			IF COUNT = "10000" THEN
				-- ZERA O CONTADOR
				COUNT := (OTHERS => '0');
			ELSE
				-- ATRIBUI O CONTADOR À SAÍDA, NO FORMATO '0000'
				S <= COUNT;
				-- INCREMENTA O CONTADOR
				COUNT := COUNT + 1;
			END IF;
			-- SE O LOAD (CARREGAR) FOR 1, ENTÃO O CONTADOR RECEBE A ENTRADA
			IF LOAD = '1' THEN
				-- ATRIBUI O DIN AO CONTADOR
				COUNT := DIN;
			END IF;
		END IF;
	END PROCESS;
END CONTADOR4BITS_ARCH;