LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY PORTA_AND IS
	PORT(
		E1: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		CLK: IN STD_LOGIC;
		S: OUT STD_LOGIC_VECTOR(7 DOWNTO 0) -- NÃO TEM ;
	);
END PORTA_AND;

ARCHITECTURE PORTA_AND_ARCH OF PORTA_AND IS
SIGNAL AUX: STD_LOGIC_VECTOR(7 DOWNTO 0);
BEGIN
	PROCESS(CLK, E1)
	BEGIN
		IF (CLK'EVENT AND CLK = '1') THEN
			AUX <= E1;
		END IF;
	END PROCESS;
	S <= AUX;
END PORTA_AND_ARCH;