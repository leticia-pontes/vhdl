LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY TB_CONTADOR4BITS IS
END TB_CONTADOR4BITS;

ARCHITECTURE TB OF TB_CONTADOR4BITS IS
	COMPONENT CONTADOR4BITS IS
	PORT(
		CLK, RST, LOAD: IN STD_LOGIC;
		DIN: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		S: OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
   END COMPONENT;
   
   SIGNAL CLK, RST, LOAD, PAUSE: STD_LOGIC;
   SIGNAL DIN, S: STD_LOGIC_VECTOR(3 DOWNTO 0);
BEGIN
	DUT: CONTADOR4BITS
	PORT MAP (CLK  => CLK,
             RST  => RST,
             LOAD => LOAD,
             DIN  => DIN,
             S    => S);
	
	CLK <= NOT CLK AFTER 50 NS WHEN PAUSE = '0' ELSE '0';
	
   STIMULI: PROCESS
   BEGIN
		PAUSE <= '0';
		
      RST  <= '0';
      LOAD <= '0';
      DIN  <= (OTHERS => '0');
		WAIT FOR 100 NS;
		
		RST <= '1';
		WAIT FOR 100 NS;
		
		RST <= '0';
		WAIT FOR 2000 NS;
     
		DIN  <= "0101";
		LOAD <= '1';
		WAIT FOR 100 NS;
      
		LOAD <= '0';
      WAIT FOR 2000 NS;
		
		PAUSE <= '1';
		WAIT;
   END PROCESS;	 
END TB;
