LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY RAM IS
	PORT(
		-- CLOCK, RESET, GRAVAÇÃO
		CLK, RST, WRITE_RAM: IN STD_LOGIC;
		-- ENDEREÇO DE DADO
		RAM_ADDR: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		-- ENTRADA DE DADO
		RAM_DATAIN: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		-- SAÍDA DE DADO
		RAM_DATAOUT: OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END RAM;

ARCHITECTURE RTL OF RAM IS
	TYPE BLOCK1_ARRAY IS ARRAY(31 DOWNTO 0) OF STD_LOGIC_VECTOR(7 DOWNTO 0); -- ARRAY PERSONALIZADO, 32 POSIÇÕES
	
	-- ARRAY BLOCK1 DO TIPO BLOCK1_ARRAY (PERSONALIZADO)
	SIGNAL BLOCK1: BLOCK1_ARRAY;
	-- INDICA A PRIMEIRA EXECUÇÃO (?)
	SIGNAL FIRST: BOOLEAN := TRUE;
BEGIN
	PROCESS(CLK, RST)
	BEGIN
		-- SE O RESET FOR ATIVADO, RESETA O "FIRST"
		IF RST = '1' THEN
			FIRST <= TRUE;
		
		-- QUANDO O CLOCK ESTIVER EM 1
		ELSIF CLK'EVENT AND CLK = '1' THEN
			-- SE "FIRST" É VERDADEIRO, QUER DIZER QUE É A PRIMEIRA EXECUÇÃO (?), LOGO O ARRAY É INICIALIZADO COM "00000000", NESSE CASO
			IF FIRST THEN
				FOR i IN 0 TO 31 LOOP
					BLOCK1(i) <= (OTHERS => '0');
				END LOOP;
				-- COLOCA O "FIRST" EM 0 PARA INDICAR QUE JÁ FOI EXECUTADO 1 VEZ
				FIRST <= FALSE;
			END IF;
			
			-- SE A GRAVAÇÃO ESTIVER EM 1
			IF WRITE_RAM = '1' THEN
				-- O ARRAY É PREENCHIDO COM A ENTRADA DE DADO (LEVA O ENDEREÇO DA MEMÓRIA COMO PARÂMETRO)
				BLOCK1(TO_INTEGER(UNSIGNED(RAM_ADDR))) <= RAM_DATAIN;
			END IF;
		END IF;
	END PROCESS;
	
	-- A SAÍDA RECEBE O ARRAY PREENCHIDO (O ARRAY LEVA O ENDEREÇO DA MEMÓRIA COMO PARÂMETRO)
	RAM_DATAOUT <= BLOCK1(TO_INTEGER(UNSIGNED(RAM_ADDR)));
END RTL;