LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY SUBTRAIR IS
	PORT (E1, E2: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			S: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END SUBTRAIR;

ARCHITECTURE SUBTRAIR_ARCH OF SUBTRAIR IS
BEGIN
	S <= E1 - E2;
END SUBTRAIR_ARCH;